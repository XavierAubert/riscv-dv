// TODO: Add custom instruction format there
// X0_FORMAT,
// X1_FORMAT,
