// TODO: Add custom instruction categories there
// MY_CUSTOM_CATEGORY_0,
// MY_CUSTOM_CATEGORY_1,
